`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/08/2021 11:45:17 PM
// Design Name: 
// Module Name: SIEMPRE4
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SIEMPRE4(
    output reg [31:0] SIEMPRE4
    );
    
    initial
        assign SIEMPRE4 = 4;
    
endmodule
